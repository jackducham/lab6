module datapath
(
	input logic GATEPC,
					GATEMDR,
					LD_MAR,
					LD_MDR,
					LD_IR,
					LD_PC,
					MIO_EN,
	input logic[1:0] PCMUX,
	input logic[15:0] MDR_In, MAR, MDR, PC, IR,
	
							
);



endmodule
